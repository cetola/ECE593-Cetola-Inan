/*
Low level (grey box) checker.
*/

module vip_checker;
//STUB
endmodule