class coverage;

    //TODO:Stub
    function new ();
    endfunction : new

    //TODO: Stub
    task execute();
    endtask : execute
endclass : coverage

