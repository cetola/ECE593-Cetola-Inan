class tester;

    virtual vip_bfm bfm;

    function new (virtual vip_bfm b);
        bfm = b;
    endfunction : new
    
    //TODO: Stub
    task execute();
    endtask : execute
endclass : tester

